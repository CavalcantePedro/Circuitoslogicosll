module lista1ex2
(input logic [7:0] entrada);



endmodule